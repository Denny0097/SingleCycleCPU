module SingleCycleCPU(
    input clk,                
    input reset               
);




endmodule