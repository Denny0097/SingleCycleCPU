module ALU (
    input   [31:0]      input1,
    input   [31:0]      input2,
    input   [3:0]       alu_controll,   // 
    output  reg [31:0]  reslut,
);
        



    
endmodule